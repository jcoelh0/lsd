library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity ROM_16_8 is
   port(address : in  std_logic_vector(3 downto 0);
        dataOut : out std_logic_vector(7 downto 0));
end ROM_16_8;

architecture RTL of ROM_16_8 is
   subtype TDataWord is std_logic_vector(7 downto 0);
   type TROM is array (0 to 15) of TDataWord;
   constant c_memory: TROM := (x"0F", x"1F", x"2F", x"3F",
                               x"AF", x"DF", x"4F", x"7F",
                               x"BF", x"EF", x"5F", x"8F",
                               x"CF", x"FF", x"6F", x"9F");

   begin
      dataOut <= c_memory(to_integer(unsigned(address)));
end RTL;